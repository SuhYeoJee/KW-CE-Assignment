`timescale 1ns/100ps

module tb_ha;
	reg a;
	reg b;
	wire s;
	wire co;
	ha ha(.a(a),.b(b),.s(s),.co(co)); // half adder
	
	initial
	begin
	a=0; b=0; //exhaustive verification
   #10; b=1;
   #10; a=1;
   #10; b=0;
   #10;
   end
endmodule
