module _4_to_23_decoder(d,q); // 4 to 23 decoder
	input [15:0] d;
	output reg [22:0] q;
	
	always@(d) begin
		if(d[15:8] == 8'h01) begin
			if(d[7:4] == 4'b0000) begin	// 9 ~ 0
				q[22:10] = 12'b0;
				case(d[3:0])
					4'b0000: q[9:0] = 10'b0000000001;
					4'b0001: q[9:0] = 10'b0000000010;
					4'b0010: q[9:0] = 10'b0000000100;
					4'b0011: q[9:0] = 10'b0000001000;
					4'b0100: q[9:0] = 10'b0000010000;
					4'b0101: q[9:0] = 10'b0000100000;
					4'b0110: q[9:0] = 10'b0001000000;
					4'b0111: q[9:0] = 10'b0010000000;
					4'b1000: q[9:0] = 10'b0100000000;
					4'b1001: q[9:0] = 10'b1000000000;
					default: q[9:0] = 10'hx;
				endcase
			end
			else if(d[7:4] == 4'b0001) begin // 19 ~ 10
				q[22:20] = 3'b0;
				q[9:0] = 10'b0;
				case(d[3:0])
					4'b0000: q[19:10] = 10'b0000000001;
					4'b0001: q[19:10] = 10'b0000000010;
					4'b0010: q[19:10] = 10'b0000000100;
					4'b0011: q[19:10] = 10'b0000001000;
					4'b0100: q[19:10] = 10'b0000010000;
					4'b0101: q[19:10] = 10'b0000100000;
					4'b0110: q[19:10] = 10'b0001000000;
					4'b0111: q[19:10] = 10'b0010000000;
					4'b1000: q[19:10] = 10'b0100000000;
					4'b1001: q[19:10] = 10'b1000000000;
					default: q[19:10] = 10'hx;
				endcase
			end
			else if(d[7:4] == 4'b0010) begin //22 ~ 20
				q[19:0] = 20'b0;
				case(d[3:0])
					4'b0000: q[22:20] = 3'b001;
					4'b0001: q[22:20] = 3'b010;
					4'b0010: q[22:20] = 3'b100;
					default: q[22:20] = 3'hx;
				endcase
			end
			else q = 23'bx;
		end
		else q = 23'bx;
	end
endmodule